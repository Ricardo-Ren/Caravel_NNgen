magic
tech sky130A
magscale 1 2
timestamp 1654153920
<< obsli1 >>
rect 1104 2159 578864 597329
<< obsm1 >>
rect 1104 2128 578864 597360
<< metal2 >>
rect 2410 599200 2466 600000
rect 7194 599200 7250 600000
rect 11978 599200 12034 600000
rect 16762 599200 16818 600000
rect 21546 599200 21602 600000
rect 26330 599200 26386 600000
rect 31114 599200 31170 600000
rect 35898 599200 35954 600000
rect 40682 599200 40738 600000
rect 45466 599200 45522 600000
rect 50250 599200 50306 600000
rect 55126 599200 55182 600000
rect 59910 599200 59966 600000
rect 64694 599200 64750 600000
rect 69478 599200 69534 600000
rect 74262 599200 74318 600000
rect 79046 599200 79102 600000
rect 83830 599200 83886 600000
rect 88614 599200 88670 600000
rect 93398 599200 93454 600000
rect 98182 599200 98238 600000
rect 103058 599200 103114 600000
rect 107842 599200 107898 600000
rect 112626 599200 112682 600000
rect 117410 599200 117466 600000
rect 122194 599200 122250 600000
rect 126978 599200 127034 600000
rect 131762 599200 131818 600000
rect 136546 599200 136602 600000
rect 141330 599200 141386 600000
rect 146114 599200 146170 600000
rect 150990 599200 151046 600000
rect 155774 599200 155830 600000
rect 160558 599200 160614 600000
rect 165342 599200 165398 600000
rect 170126 599200 170182 600000
rect 174910 599200 174966 600000
rect 179694 599200 179750 600000
rect 184478 599200 184534 600000
rect 189262 599200 189318 600000
rect 194046 599200 194102 600000
rect 198922 599200 198978 600000
rect 203706 599200 203762 600000
rect 208490 599200 208546 600000
rect 213274 599200 213330 600000
rect 218058 599200 218114 600000
rect 222842 599200 222898 600000
rect 227626 599200 227682 600000
rect 232410 599200 232466 600000
rect 237194 599200 237250 600000
rect 241978 599200 242034 600000
rect 246854 599200 246910 600000
rect 251638 599200 251694 600000
rect 256422 599200 256478 600000
rect 261206 599200 261262 600000
rect 265990 599200 266046 600000
rect 270774 599200 270830 600000
rect 275558 599200 275614 600000
rect 280342 599200 280398 600000
rect 285126 599200 285182 600000
rect 289910 599200 289966 600000
rect 294786 599200 294842 600000
rect 299570 599200 299626 600000
rect 304354 599200 304410 600000
rect 309138 599200 309194 600000
rect 313922 599200 313978 600000
rect 318706 599200 318762 600000
rect 323490 599200 323546 600000
rect 328274 599200 328330 600000
rect 333058 599200 333114 600000
rect 337842 599200 337898 600000
rect 342718 599200 342774 600000
rect 347502 599200 347558 600000
rect 352286 599200 352342 600000
rect 357070 599200 357126 600000
rect 361854 599200 361910 600000
rect 366638 599200 366694 600000
rect 371422 599200 371478 600000
rect 376206 599200 376262 600000
rect 380990 599200 381046 600000
rect 385774 599200 385830 600000
rect 390650 599200 390706 600000
rect 395434 599200 395490 600000
rect 400218 599200 400274 600000
rect 405002 599200 405058 600000
rect 409786 599200 409842 600000
rect 414570 599200 414626 600000
rect 419354 599200 419410 600000
rect 424138 599200 424194 600000
rect 428922 599200 428978 600000
rect 433706 599200 433762 600000
rect 438582 599200 438638 600000
rect 443366 599200 443422 600000
rect 448150 599200 448206 600000
rect 452934 599200 452990 600000
rect 457718 599200 457774 600000
rect 462502 599200 462558 600000
rect 467286 599200 467342 600000
rect 472070 599200 472126 600000
rect 476854 599200 476910 600000
rect 481638 599200 481694 600000
rect 486514 599200 486570 600000
rect 491298 599200 491354 600000
rect 496082 599200 496138 600000
rect 500866 599200 500922 600000
rect 505650 599200 505706 600000
rect 510434 599200 510490 600000
rect 515218 599200 515274 600000
rect 520002 599200 520058 600000
rect 524786 599200 524842 600000
rect 529570 599200 529626 600000
rect 534446 599200 534502 600000
rect 539230 599200 539286 600000
rect 544014 599200 544070 600000
rect 548798 599200 548854 600000
rect 553582 599200 553638 600000
rect 558366 599200 558422 600000
rect 563150 599200 563206 600000
rect 567934 599200 567990 600000
rect 572718 599200 572774 600000
rect 577502 599200 577558 600000
rect 570 0 626 800
rect 1674 0 1730 800
rect 2870 0 2926 800
rect 4066 0 4122 800
rect 5170 0 5226 800
rect 6366 0 6422 800
rect 7562 0 7618 800
rect 8666 0 8722 800
rect 9862 0 9918 800
rect 11058 0 11114 800
rect 12162 0 12218 800
rect 13358 0 13414 800
rect 14554 0 14610 800
rect 15658 0 15714 800
rect 16854 0 16910 800
rect 18050 0 18106 800
rect 19154 0 19210 800
rect 20350 0 20406 800
rect 21546 0 21602 800
rect 22650 0 22706 800
rect 23846 0 23902 800
rect 25042 0 25098 800
rect 26238 0 26294 800
rect 27342 0 27398 800
rect 28538 0 28594 800
rect 29734 0 29790 800
rect 30838 0 30894 800
rect 32034 0 32090 800
rect 33230 0 33286 800
rect 34334 0 34390 800
rect 35530 0 35586 800
rect 36726 0 36782 800
rect 37830 0 37886 800
rect 39026 0 39082 800
rect 40222 0 40278 800
rect 41326 0 41382 800
rect 42522 0 42578 800
rect 43718 0 43774 800
rect 44822 0 44878 800
rect 46018 0 46074 800
rect 47214 0 47270 800
rect 48410 0 48466 800
rect 49514 0 49570 800
rect 50710 0 50766 800
rect 51906 0 51962 800
rect 53010 0 53066 800
rect 54206 0 54262 800
rect 55402 0 55458 800
rect 56506 0 56562 800
rect 57702 0 57758 800
rect 58898 0 58954 800
rect 60002 0 60058 800
rect 61198 0 61254 800
rect 62394 0 62450 800
rect 63498 0 63554 800
rect 64694 0 64750 800
rect 65890 0 65946 800
rect 66994 0 67050 800
rect 68190 0 68246 800
rect 69386 0 69442 800
rect 70582 0 70638 800
rect 71686 0 71742 800
rect 72882 0 72938 800
rect 74078 0 74134 800
rect 75182 0 75238 800
rect 76378 0 76434 800
rect 77574 0 77630 800
rect 78678 0 78734 800
rect 79874 0 79930 800
rect 81070 0 81126 800
rect 82174 0 82230 800
rect 83370 0 83426 800
rect 84566 0 84622 800
rect 85670 0 85726 800
rect 86866 0 86922 800
rect 88062 0 88118 800
rect 89166 0 89222 800
rect 90362 0 90418 800
rect 91558 0 91614 800
rect 92754 0 92810 800
rect 93858 0 93914 800
rect 95054 0 95110 800
rect 96250 0 96306 800
rect 97354 0 97410 800
rect 98550 0 98606 800
rect 99746 0 99802 800
rect 100850 0 100906 800
rect 102046 0 102102 800
rect 103242 0 103298 800
rect 104346 0 104402 800
rect 105542 0 105598 800
rect 106738 0 106794 800
rect 107842 0 107898 800
rect 109038 0 109094 800
rect 110234 0 110290 800
rect 111338 0 111394 800
rect 112534 0 112590 800
rect 113730 0 113786 800
rect 114926 0 114982 800
rect 116030 0 116086 800
rect 117226 0 117282 800
rect 118422 0 118478 800
rect 119526 0 119582 800
rect 120722 0 120778 800
rect 121918 0 121974 800
rect 123022 0 123078 800
rect 124218 0 124274 800
rect 125414 0 125470 800
rect 126518 0 126574 800
rect 127714 0 127770 800
rect 128910 0 128966 800
rect 130014 0 130070 800
rect 131210 0 131266 800
rect 132406 0 132462 800
rect 133510 0 133566 800
rect 134706 0 134762 800
rect 135902 0 135958 800
rect 137098 0 137154 800
rect 138202 0 138258 800
rect 139398 0 139454 800
rect 140594 0 140650 800
rect 141698 0 141754 800
rect 142894 0 142950 800
rect 144090 0 144146 800
rect 145194 0 145250 800
rect 146390 0 146446 800
rect 147586 0 147642 800
rect 148690 0 148746 800
rect 149886 0 149942 800
rect 151082 0 151138 800
rect 152186 0 152242 800
rect 153382 0 153438 800
rect 154578 0 154634 800
rect 155682 0 155738 800
rect 156878 0 156934 800
rect 158074 0 158130 800
rect 159270 0 159326 800
rect 160374 0 160430 800
rect 161570 0 161626 800
rect 162766 0 162822 800
rect 163870 0 163926 800
rect 165066 0 165122 800
rect 166262 0 166318 800
rect 167366 0 167422 800
rect 168562 0 168618 800
rect 169758 0 169814 800
rect 170862 0 170918 800
rect 172058 0 172114 800
rect 173254 0 173310 800
rect 174358 0 174414 800
rect 175554 0 175610 800
rect 176750 0 176806 800
rect 177854 0 177910 800
rect 179050 0 179106 800
rect 180246 0 180302 800
rect 181442 0 181498 800
rect 182546 0 182602 800
rect 183742 0 183798 800
rect 184938 0 184994 800
rect 186042 0 186098 800
rect 187238 0 187294 800
rect 188434 0 188490 800
rect 189538 0 189594 800
rect 190734 0 190790 800
rect 191930 0 191986 800
rect 193034 0 193090 800
rect 194230 0 194286 800
rect 195426 0 195482 800
rect 196530 0 196586 800
rect 197726 0 197782 800
rect 198922 0 198978 800
rect 200026 0 200082 800
rect 201222 0 201278 800
rect 202418 0 202474 800
rect 203614 0 203670 800
rect 204718 0 204774 800
rect 205914 0 205970 800
rect 207110 0 207166 800
rect 208214 0 208270 800
rect 209410 0 209466 800
rect 210606 0 210662 800
rect 211710 0 211766 800
rect 212906 0 212962 800
rect 214102 0 214158 800
rect 215206 0 215262 800
rect 216402 0 216458 800
rect 217598 0 217654 800
rect 218702 0 218758 800
rect 219898 0 219954 800
rect 221094 0 221150 800
rect 222198 0 222254 800
rect 223394 0 223450 800
rect 224590 0 224646 800
rect 225786 0 225842 800
rect 226890 0 226946 800
rect 228086 0 228142 800
rect 229282 0 229338 800
rect 230386 0 230442 800
rect 231582 0 231638 800
rect 232778 0 232834 800
rect 233882 0 233938 800
rect 235078 0 235134 800
rect 236274 0 236330 800
rect 237378 0 237434 800
rect 238574 0 238630 800
rect 239770 0 239826 800
rect 240874 0 240930 800
rect 242070 0 242126 800
rect 243266 0 243322 800
rect 244370 0 244426 800
rect 245566 0 245622 800
rect 246762 0 246818 800
rect 247958 0 248014 800
rect 249062 0 249118 800
rect 250258 0 250314 800
rect 251454 0 251510 800
rect 252558 0 252614 800
rect 253754 0 253810 800
rect 254950 0 255006 800
rect 256054 0 256110 800
rect 257250 0 257306 800
rect 258446 0 258502 800
rect 259550 0 259606 800
rect 260746 0 260802 800
rect 261942 0 261998 800
rect 263046 0 263102 800
rect 264242 0 264298 800
rect 265438 0 265494 800
rect 266542 0 266598 800
rect 267738 0 267794 800
rect 268934 0 268990 800
rect 270130 0 270186 800
rect 271234 0 271290 800
rect 272430 0 272486 800
rect 273626 0 273682 800
rect 274730 0 274786 800
rect 275926 0 275982 800
rect 277122 0 277178 800
rect 278226 0 278282 800
rect 279422 0 279478 800
rect 280618 0 280674 800
rect 281722 0 281778 800
rect 282918 0 282974 800
rect 284114 0 284170 800
rect 285218 0 285274 800
rect 286414 0 286470 800
rect 287610 0 287666 800
rect 288714 0 288770 800
rect 289910 0 289966 800
rect 291106 0 291162 800
rect 292302 0 292358 800
rect 293406 0 293462 800
rect 294602 0 294658 800
rect 295798 0 295854 800
rect 296902 0 296958 800
rect 298098 0 298154 800
rect 299294 0 299350 800
rect 300398 0 300454 800
rect 301594 0 301650 800
rect 302790 0 302846 800
rect 303894 0 303950 800
rect 305090 0 305146 800
rect 306286 0 306342 800
rect 307390 0 307446 800
rect 308586 0 308642 800
rect 309782 0 309838 800
rect 310886 0 310942 800
rect 312082 0 312138 800
rect 313278 0 313334 800
rect 314474 0 314530 800
rect 315578 0 315634 800
rect 316774 0 316830 800
rect 317970 0 318026 800
rect 319074 0 319130 800
rect 320270 0 320326 800
rect 321466 0 321522 800
rect 322570 0 322626 800
rect 323766 0 323822 800
rect 324962 0 325018 800
rect 326066 0 326122 800
rect 327262 0 327318 800
rect 328458 0 328514 800
rect 329562 0 329618 800
rect 330758 0 330814 800
rect 331954 0 332010 800
rect 333058 0 333114 800
rect 334254 0 334310 800
rect 335450 0 335506 800
rect 336646 0 336702 800
rect 337750 0 337806 800
rect 338946 0 339002 800
rect 340142 0 340198 800
rect 341246 0 341302 800
rect 342442 0 342498 800
rect 343638 0 343694 800
rect 344742 0 344798 800
rect 345938 0 345994 800
rect 347134 0 347190 800
rect 348238 0 348294 800
rect 349434 0 349490 800
rect 350630 0 350686 800
rect 351734 0 351790 800
rect 352930 0 352986 800
rect 354126 0 354182 800
rect 355230 0 355286 800
rect 356426 0 356482 800
rect 357622 0 357678 800
rect 358818 0 358874 800
rect 359922 0 359978 800
rect 361118 0 361174 800
rect 362314 0 362370 800
rect 363418 0 363474 800
rect 364614 0 364670 800
rect 365810 0 365866 800
rect 366914 0 366970 800
rect 368110 0 368166 800
rect 369306 0 369362 800
rect 370410 0 370466 800
rect 371606 0 371662 800
rect 372802 0 372858 800
rect 373906 0 373962 800
rect 375102 0 375158 800
rect 376298 0 376354 800
rect 377402 0 377458 800
rect 378598 0 378654 800
rect 379794 0 379850 800
rect 380990 0 381046 800
rect 382094 0 382150 800
rect 383290 0 383346 800
rect 384486 0 384542 800
rect 385590 0 385646 800
rect 386786 0 386842 800
rect 387982 0 388038 800
rect 389086 0 389142 800
rect 390282 0 390338 800
rect 391478 0 391534 800
rect 392582 0 392638 800
rect 393778 0 393834 800
rect 394974 0 395030 800
rect 396078 0 396134 800
rect 397274 0 397330 800
rect 398470 0 398526 800
rect 399574 0 399630 800
rect 400770 0 400826 800
rect 401966 0 402022 800
rect 403162 0 403218 800
rect 404266 0 404322 800
rect 405462 0 405518 800
rect 406658 0 406714 800
rect 407762 0 407818 800
rect 408958 0 409014 800
rect 410154 0 410210 800
rect 411258 0 411314 800
rect 412454 0 412510 800
rect 413650 0 413706 800
rect 414754 0 414810 800
rect 415950 0 416006 800
rect 417146 0 417202 800
rect 418250 0 418306 800
rect 419446 0 419502 800
rect 420642 0 420698 800
rect 421746 0 421802 800
rect 422942 0 422998 800
rect 424138 0 424194 800
rect 425334 0 425390 800
rect 426438 0 426494 800
rect 427634 0 427690 800
rect 428830 0 428886 800
rect 429934 0 429990 800
rect 431130 0 431186 800
rect 432326 0 432382 800
rect 433430 0 433486 800
rect 434626 0 434682 800
rect 435822 0 435878 800
rect 436926 0 436982 800
rect 438122 0 438178 800
rect 439318 0 439374 800
rect 440422 0 440478 800
rect 441618 0 441674 800
rect 442814 0 442870 800
rect 443918 0 443974 800
rect 445114 0 445170 800
rect 446310 0 446366 800
rect 447506 0 447562 800
rect 448610 0 448666 800
rect 449806 0 449862 800
rect 451002 0 451058 800
rect 452106 0 452162 800
rect 453302 0 453358 800
rect 454498 0 454554 800
rect 455602 0 455658 800
rect 456798 0 456854 800
rect 457994 0 458050 800
rect 459098 0 459154 800
rect 460294 0 460350 800
rect 461490 0 461546 800
rect 462594 0 462650 800
rect 463790 0 463846 800
rect 464986 0 465042 800
rect 466090 0 466146 800
rect 467286 0 467342 800
rect 468482 0 468538 800
rect 469678 0 469734 800
rect 470782 0 470838 800
rect 471978 0 472034 800
rect 473174 0 473230 800
rect 474278 0 474334 800
rect 475474 0 475530 800
rect 476670 0 476726 800
rect 477774 0 477830 800
rect 478970 0 479026 800
rect 480166 0 480222 800
rect 481270 0 481326 800
rect 482466 0 482522 800
rect 483662 0 483718 800
rect 484766 0 484822 800
rect 485962 0 486018 800
rect 487158 0 487214 800
rect 488262 0 488318 800
rect 489458 0 489514 800
rect 490654 0 490710 800
rect 491850 0 491906 800
rect 492954 0 493010 800
rect 494150 0 494206 800
rect 495346 0 495402 800
rect 496450 0 496506 800
rect 497646 0 497702 800
rect 498842 0 498898 800
rect 499946 0 500002 800
rect 501142 0 501198 800
rect 502338 0 502394 800
rect 503442 0 503498 800
rect 504638 0 504694 800
rect 505834 0 505890 800
rect 506938 0 506994 800
rect 508134 0 508190 800
rect 509330 0 509386 800
rect 510434 0 510490 800
rect 511630 0 511686 800
rect 512826 0 512882 800
rect 514022 0 514078 800
rect 515126 0 515182 800
rect 516322 0 516378 800
rect 517518 0 517574 800
rect 518622 0 518678 800
rect 519818 0 519874 800
rect 521014 0 521070 800
rect 522118 0 522174 800
rect 523314 0 523370 800
rect 524510 0 524566 800
rect 525614 0 525670 800
rect 526810 0 526866 800
rect 528006 0 528062 800
rect 529110 0 529166 800
rect 530306 0 530362 800
rect 531502 0 531558 800
rect 532606 0 532662 800
rect 533802 0 533858 800
rect 534998 0 535054 800
rect 536194 0 536250 800
rect 537298 0 537354 800
rect 538494 0 538550 800
rect 539690 0 539746 800
rect 540794 0 540850 800
rect 541990 0 542046 800
rect 543186 0 543242 800
rect 544290 0 544346 800
rect 545486 0 545542 800
rect 546682 0 546738 800
rect 547786 0 547842 800
rect 548982 0 549038 800
rect 550178 0 550234 800
rect 551282 0 551338 800
rect 552478 0 552534 800
rect 553674 0 553730 800
rect 554778 0 554834 800
rect 555974 0 556030 800
rect 557170 0 557226 800
rect 558366 0 558422 800
rect 559470 0 559526 800
rect 560666 0 560722 800
rect 561862 0 561918 800
rect 562966 0 563022 800
rect 564162 0 564218 800
rect 565358 0 565414 800
rect 566462 0 566518 800
rect 567658 0 567714 800
rect 568854 0 568910 800
rect 569958 0 570014 800
rect 571154 0 571210 800
rect 572350 0 572406 800
rect 573454 0 573510 800
rect 574650 0 574706 800
rect 575846 0 575902 800
rect 576950 0 577006 800
rect 578146 0 578202 800
rect 579342 0 579398 800
<< obsm2 >>
rect 570 599144 2354 599298
rect 2522 599144 7138 599298
rect 7306 599144 11922 599298
rect 12090 599144 16706 599298
rect 16874 599144 21490 599298
rect 21658 599144 26274 599298
rect 26442 599144 31058 599298
rect 31226 599144 35842 599298
rect 36010 599144 40626 599298
rect 40794 599144 45410 599298
rect 45578 599144 50194 599298
rect 50362 599144 55070 599298
rect 55238 599144 59854 599298
rect 60022 599144 64638 599298
rect 64806 599144 69422 599298
rect 69590 599144 74206 599298
rect 74374 599144 78990 599298
rect 79158 599144 83774 599298
rect 83942 599144 88558 599298
rect 88726 599144 93342 599298
rect 93510 599144 98126 599298
rect 98294 599144 103002 599298
rect 103170 599144 107786 599298
rect 107954 599144 112570 599298
rect 112738 599144 117354 599298
rect 117522 599144 122138 599298
rect 122306 599144 126922 599298
rect 127090 599144 131706 599298
rect 131874 599144 136490 599298
rect 136658 599144 141274 599298
rect 141442 599144 146058 599298
rect 146226 599144 150934 599298
rect 151102 599144 155718 599298
rect 155886 599144 160502 599298
rect 160670 599144 165286 599298
rect 165454 599144 170070 599298
rect 170238 599144 174854 599298
rect 175022 599144 179638 599298
rect 179806 599144 184422 599298
rect 184590 599144 189206 599298
rect 189374 599144 193990 599298
rect 194158 599144 198866 599298
rect 199034 599144 203650 599298
rect 203818 599144 208434 599298
rect 208602 599144 213218 599298
rect 213386 599144 218002 599298
rect 218170 599144 222786 599298
rect 222954 599144 227570 599298
rect 227738 599144 232354 599298
rect 232522 599144 237138 599298
rect 237306 599144 241922 599298
rect 242090 599144 246798 599298
rect 246966 599144 251582 599298
rect 251750 599144 256366 599298
rect 256534 599144 261150 599298
rect 261318 599144 265934 599298
rect 266102 599144 270718 599298
rect 270886 599144 275502 599298
rect 275670 599144 280286 599298
rect 280454 599144 285070 599298
rect 285238 599144 289854 599298
rect 290022 599144 294730 599298
rect 294898 599144 299514 599298
rect 299682 599144 304298 599298
rect 304466 599144 309082 599298
rect 309250 599144 313866 599298
rect 314034 599144 318650 599298
rect 318818 599144 323434 599298
rect 323602 599144 328218 599298
rect 328386 599144 333002 599298
rect 333170 599144 337786 599298
rect 337954 599144 342662 599298
rect 342830 599144 347446 599298
rect 347614 599144 352230 599298
rect 352398 599144 357014 599298
rect 357182 599144 361798 599298
rect 361966 599144 366582 599298
rect 366750 599144 371366 599298
rect 371534 599144 376150 599298
rect 376318 599144 380934 599298
rect 381102 599144 385718 599298
rect 385886 599144 390594 599298
rect 390762 599144 395378 599298
rect 395546 599144 400162 599298
rect 400330 599144 404946 599298
rect 405114 599144 409730 599298
rect 409898 599144 414514 599298
rect 414682 599144 419298 599298
rect 419466 599144 424082 599298
rect 424250 599144 428866 599298
rect 429034 599144 433650 599298
rect 433818 599144 438526 599298
rect 438694 599144 443310 599298
rect 443478 599144 448094 599298
rect 448262 599144 452878 599298
rect 453046 599144 457662 599298
rect 457830 599144 462446 599298
rect 462614 599144 467230 599298
rect 467398 599144 472014 599298
rect 472182 599144 476798 599298
rect 476966 599144 481582 599298
rect 481750 599144 486458 599298
rect 486626 599144 491242 599298
rect 491410 599144 496026 599298
rect 496194 599144 500810 599298
rect 500978 599144 505594 599298
rect 505762 599144 510378 599298
rect 510546 599144 515162 599298
rect 515330 599144 519946 599298
rect 520114 599144 524730 599298
rect 524898 599144 529514 599298
rect 529682 599144 534390 599298
rect 534558 599144 539174 599298
rect 539342 599144 543958 599298
rect 544126 599144 548742 599298
rect 548910 599144 553526 599298
rect 553694 599144 558310 599298
rect 558478 599144 563094 599298
rect 563262 599144 567878 599298
rect 568046 599144 572662 599298
rect 572830 599144 577446 599298
rect 577614 599144 577742 599298
rect 570 856 577742 599144
rect 682 800 1618 856
rect 1786 800 2814 856
rect 2982 800 4010 856
rect 4178 800 5114 856
rect 5282 800 6310 856
rect 6478 800 7506 856
rect 7674 800 8610 856
rect 8778 800 9806 856
rect 9974 800 11002 856
rect 11170 800 12106 856
rect 12274 800 13302 856
rect 13470 800 14498 856
rect 14666 800 15602 856
rect 15770 800 16798 856
rect 16966 800 17994 856
rect 18162 800 19098 856
rect 19266 800 20294 856
rect 20462 800 21490 856
rect 21658 800 22594 856
rect 22762 800 23790 856
rect 23958 800 24986 856
rect 25154 800 26182 856
rect 26350 800 27286 856
rect 27454 800 28482 856
rect 28650 800 29678 856
rect 29846 800 30782 856
rect 30950 800 31978 856
rect 32146 800 33174 856
rect 33342 800 34278 856
rect 34446 800 35474 856
rect 35642 800 36670 856
rect 36838 800 37774 856
rect 37942 800 38970 856
rect 39138 800 40166 856
rect 40334 800 41270 856
rect 41438 800 42466 856
rect 42634 800 43662 856
rect 43830 800 44766 856
rect 44934 800 45962 856
rect 46130 800 47158 856
rect 47326 800 48354 856
rect 48522 800 49458 856
rect 49626 800 50654 856
rect 50822 800 51850 856
rect 52018 800 52954 856
rect 53122 800 54150 856
rect 54318 800 55346 856
rect 55514 800 56450 856
rect 56618 800 57646 856
rect 57814 800 58842 856
rect 59010 800 59946 856
rect 60114 800 61142 856
rect 61310 800 62338 856
rect 62506 800 63442 856
rect 63610 800 64638 856
rect 64806 800 65834 856
rect 66002 800 66938 856
rect 67106 800 68134 856
rect 68302 800 69330 856
rect 69498 800 70526 856
rect 70694 800 71630 856
rect 71798 800 72826 856
rect 72994 800 74022 856
rect 74190 800 75126 856
rect 75294 800 76322 856
rect 76490 800 77518 856
rect 77686 800 78622 856
rect 78790 800 79818 856
rect 79986 800 81014 856
rect 81182 800 82118 856
rect 82286 800 83314 856
rect 83482 800 84510 856
rect 84678 800 85614 856
rect 85782 800 86810 856
rect 86978 800 88006 856
rect 88174 800 89110 856
rect 89278 800 90306 856
rect 90474 800 91502 856
rect 91670 800 92698 856
rect 92866 800 93802 856
rect 93970 800 94998 856
rect 95166 800 96194 856
rect 96362 800 97298 856
rect 97466 800 98494 856
rect 98662 800 99690 856
rect 99858 800 100794 856
rect 100962 800 101990 856
rect 102158 800 103186 856
rect 103354 800 104290 856
rect 104458 800 105486 856
rect 105654 800 106682 856
rect 106850 800 107786 856
rect 107954 800 108982 856
rect 109150 800 110178 856
rect 110346 800 111282 856
rect 111450 800 112478 856
rect 112646 800 113674 856
rect 113842 800 114870 856
rect 115038 800 115974 856
rect 116142 800 117170 856
rect 117338 800 118366 856
rect 118534 800 119470 856
rect 119638 800 120666 856
rect 120834 800 121862 856
rect 122030 800 122966 856
rect 123134 800 124162 856
rect 124330 800 125358 856
rect 125526 800 126462 856
rect 126630 800 127658 856
rect 127826 800 128854 856
rect 129022 800 129958 856
rect 130126 800 131154 856
rect 131322 800 132350 856
rect 132518 800 133454 856
rect 133622 800 134650 856
rect 134818 800 135846 856
rect 136014 800 137042 856
rect 137210 800 138146 856
rect 138314 800 139342 856
rect 139510 800 140538 856
rect 140706 800 141642 856
rect 141810 800 142838 856
rect 143006 800 144034 856
rect 144202 800 145138 856
rect 145306 800 146334 856
rect 146502 800 147530 856
rect 147698 800 148634 856
rect 148802 800 149830 856
rect 149998 800 151026 856
rect 151194 800 152130 856
rect 152298 800 153326 856
rect 153494 800 154522 856
rect 154690 800 155626 856
rect 155794 800 156822 856
rect 156990 800 158018 856
rect 158186 800 159214 856
rect 159382 800 160318 856
rect 160486 800 161514 856
rect 161682 800 162710 856
rect 162878 800 163814 856
rect 163982 800 165010 856
rect 165178 800 166206 856
rect 166374 800 167310 856
rect 167478 800 168506 856
rect 168674 800 169702 856
rect 169870 800 170806 856
rect 170974 800 172002 856
rect 172170 800 173198 856
rect 173366 800 174302 856
rect 174470 800 175498 856
rect 175666 800 176694 856
rect 176862 800 177798 856
rect 177966 800 178994 856
rect 179162 800 180190 856
rect 180358 800 181386 856
rect 181554 800 182490 856
rect 182658 800 183686 856
rect 183854 800 184882 856
rect 185050 800 185986 856
rect 186154 800 187182 856
rect 187350 800 188378 856
rect 188546 800 189482 856
rect 189650 800 190678 856
rect 190846 800 191874 856
rect 192042 800 192978 856
rect 193146 800 194174 856
rect 194342 800 195370 856
rect 195538 800 196474 856
rect 196642 800 197670 856
rect 197838 800 198866 856
rect 199034 800 199970 856
rect 200138 800 201166 856
rect 201334 800 202362 856
rect 202530 800 203558 856
rect 203726 800 204662 856
rect 204830 800 205858 856
rect 206026 800 207054 856
rect 207222 800 208158 856
rect 208326 800 209354 856
rect 209522 800 210550 856
rect 210718 800 211654 856
rect 211822 800 212850 856
rect 213018 800 214046 856
rect 214214 800 215150 856
rect 215318 800 216346 856
rect 216514 800 217542 856
rect 217710 800 218646 856
rect 218814 800 219842 856
rect 220010 800 221038 856
rect 221206 800 222142 856
rect 222310 800 223338 856
rect 223506 800 224534 856
rect 224702 800 225730 856
rect 225898 800 226834 856
rect 227002 800 228030 856
rect 228198 800 229226 856
rect 229394 800 230330 856
rect 230498 800 231526 856
rect 231694 800 232722 856
rect 232890 800 233826 856
rect 233994 800 235022 856
rect 235190 800 236218 856
rect 236386 800 237322 856
rect 237490 800 238518 856
rect 238686 800 239714 856
rect 239882 800 240818 856
rect 240986 800 242014 856
rect 242182 800 243210 856
rect 243378 800 244314 856
rect 244482 800 245510 856
rect 245678 800 246706 856
rect 246874 800 247902 856
rect 248070 800 249006 856
rect 249174 800 250202 856
rect 250370 800 251398 856
rect 251566 800 252502 856
rect 252670 800 253698 856
rect 253866 800 254894 856
rect 255062 800 255998 856
rect 256166 800 257194 856
rect 257362 800 258390 856
rect 258558 800 259494 856
rect 259662 800 260690 856
rect 260858 800 261886 856
rect 262054 800 262990 856
rect 263158 800 264186 856
rect 264354 800 265382 856
rect 265550 800 266486 856
rect 266654 800 267682 856
rect 267850 800 268878 856
rect 269046 800 270074 856
rect 270242 800 271178 856
rect 271346 800 272374 856
rect 272542 800 273570 856
rect 273738 800 274674 856
rect 274842 800 275870 856
rect 276038 800 277066 856
rect 277234 800 278170 856
rect 278338 800 279366 856
rect 279534 800 280562 856
rect 280730 800 281666 856
rect 281834 800 282862 856
rect 283030 800 284058 856
rect 284226 800 285162 856
rect 285330 800 286358 856
rect 286526 800 287554 856
rect 287722 800 288658 856
rect 288826 800 289854 856
rect 290022 800 291050 856
rect 291218 800 292246 856
rect 292414 800 293350 856
rect 293518 800 294546 856
rect 294714 800 295742 856
rect 295910 800 296846 856
rect 297014 800 298042 856
rect 298210 800 299238 856
rect 299406 800 300342 856
rect 300510 800 301538 856
rect 301706 800 302734 856
rect 302902 800 303838 856
rect 304006 800 305034 856
rect 305202 800 306230 856
rect 306398 800 307334 856
rect 307502 800 308530 856
rect 308698 800 309726 856
rect 309894 800 310830 856
rect 310998 800 312026 856
rect 312194 800 313222 856
rect 313390 800 314418 856
rect 314586 800 315522 856
rect 315690 800 316718 856
rect 316886 800 317914 856
rect 318082 800 319018 856
rect 319186 800 320214 856
rect 320382 800 321410 856
rect 321578 800 322514 856
rect 322682 800 323710 856
rect 323878 800 324906 856
rect 325074 800 326010 856
rect 326178 800 327206 856
rect 327374 800 328402 856
rect 328570 800 329506 856
rect 329674 800 330702 856
rect 330870 800 331898 856
rect 332066 800 333002 856
rect 333170 800 334198 856
rect 334366 800 335394 856
rect 335562 800 336590 856
rect 336758 800 337694 856
rect 337862 800 338890 856
rect 339058 800 340086 856
rect 340254 800 341190 856
rect 341358 800 342386 856
rect 342554 800 343582 856
rect 343750 800 344686 856
rect 344854 800 345882 856
rect 346050 800 347078 856
rect 347246 800 348182 856
rect 348350 800 349378 856
rect 349546 800 350574 856
rect 350742 800 351678 856
rect 351846 800 352874 856
rect 353042 800 354070 856
rect 354238 800 355174 856
rect 355342 800 356370 856
rect 356538 800 357566 856
rect 357734 800 358762 856
rect 358930 800 359866 856
rect 360034 800 361062 856
rect 361230 800 362258 856
rect 362426 800 363362 856
rect 363530 800 364558 856
rect 364726 800 365754 856
rect 365922 800 366858 856
rect 367026 800 368054 856
rect 368222 800 369250 856
rect 369418 800 370354 856
rect 370522 800 371550 856
rect 371718 800 372746 856
rect 372914 800 373850 856
rect 374018 800 375046 856
rect 375214 800 376242 856
rect 376410 800 377346 856
rect 377514 800 378542 856
rect 378710 800 379738 856
rect 379906 800 380934 856
rect 381102 800 382038 856
rect 382206 800 383234 856
rect 383402 800 384430 856
rect 384598 800 385534 856
rect 385702 800 386730 856
rect 386898 800 387926 856
rect 388094 800 389030 856
rect 389198 800 390226 856
rect 390394 800 391422 856
rect 391590 800 392526 856
rect 392694 800 393722 856
rect 393890 800 394918 856
rect 395086 800 396022 856
rect 396190 800 397218 856
rect 397386 800 398414 856
rect 398582 800 399518 856
rect 399686 800 400714 856
rect 400882 800 401910 856
rect 402078 800 403106 856
rect 403274 800 404210 856
rect 404378 800 405406 856
rect 405574 800 406602 856
rect 406770 800 407706 856
rect 407874 800 408902 856
rect 409070 800 410098 856
rect 410266 800 411202 856
rect 411370 800 412398 856
rect 412566 800 413594 856
rect 413762 800 414698 856
rect 414866 800 415894 856
rect 416062 800 417090 856
rect 417258 800 418194 856
rect 418362 800 419390 856
rect 419558 800 420586 856
rect 420754 800 421690 856
rect 421858 800 422886 856
rect 423054 800 424082 856
rect 424250 800 425278 856
rect 425446 800 426382 856
rect 426550 800 427578 856
rect 427746 800 428774 856
rect 428942 800 429878 856
rect 430046 800 431074 856
rect 431242 800 432270 856
rect 432438 800 433374 856
rect 433542 800 434570 856
rect 434738 800 435766 856
rect 435934 800 436870 856
rect 437038 800 438066 856
rect 438234 800 439262 856
rect 439430 800 440366 856
rect 440534 800 441562 856
rect 441730 800 442758 856
rect 442926 800 443862 856
rect 444030 800 445058 856
rect 445226 800 446254 856
rect 446422 800 447450 856
rect 447618 800 448554 856
rect 448722 800 449750 856
rect 449918 800 450946 856
rect 451114 800 452050 856
rect 452218 800 453246 856
rect 453414 800 454442 856
rect 454610 800 455546 856
rect 455714 800 456742 856
rect 456910 800 457938 856
rect 458106 800 459042 856
rect 459210 800 460238 856
rect 460406 800 461434 856
rect 461602 800 462538 856
rect 462706 800 463734 856
rect 463902 800 464930 856
rect 465098 800 466034 856
rect 466202 800 467230 856
rect 467398 800 468426 856
rect 468594 800 469622 856
rect 469790 800 470726 856
rect 470894 800 471922 856
rect 472090 800 473118 856
rect 473286 800 474222 856
rect 474390 800 475418 856
rect 475586 800 476614 856
rect 476782 800 477718 856
rect 477886 800 478914 856
rect 479082 800 480110 856
rect 480278 800 481214 856
rect 481382 800 482410 856
rect 482578 800 483606 856
rect 483774 800 484710 856
rect 484878 800 485906 856
rect 486074 800 487102 856
rect 487270 800 488206 856
rect 488374 800 489402 856
rect 489570 800 490598 856
rect 490766 800 491794 856
rect 491962 800 492898 856
rect 493066 800 494094 856
rect 494262 800 495290 856
rect 495458 800 496394 856
rect 496562 800 497590 856
rect 497758 800 498786 856
rect 498954 800 499890 856
rect 500058 800 501086 856
rect 501254 800 502282 856
rect 502450 800 503386 856
rect 503554 800 504582 856
rect 504750 800 505778 856
rect 505946 800 506882 856
rect 507050 800 508078 856
rect 508246 800 509274 856
rect 509442 800 510378 856
rect 510546 800 511574 856
rect 511742 800 512770 856
rect 512938 800 513966 856
rect 514134 800 515070 856
rect 515238 800 516266 856
rect 516434 800 517462 856
rect 517630 800 518566 856
rect 518734 800 519762 856
rect 519930 800 520958 856
rect 521126 800 522062 856
rect 522230 800 523258 856
rect 523426 800 524454 856
rect 524622 800 525558 856
rect 525726 800 526754 856
rect 526922 800 527950 856
rect 528118 800 529054 856
rect 529222 800 530250 856
rect 530418 800 531446 856
rect 531614 800 532550 856
rect 532718 800 533746 856
rect 533914 800 534942 856
rect 535110 800 536138 856
rect 536306 800 537242 856
rect 537410 800 538438 856
rect 538606 800 539634 856
rect 539802 800 540738 856
rect 540906 800 541934 856
rect 542102 800 543130 856
rect 543298 800 544234 856
rect 544402 800 545430 856
rect 545598 800 546626 856
rect 546794 800 547730 856
rect 547898 800 548926 856
rect 549094 800 550122 856
rect 550290 800 551226 856
rect 551394 800 552422 856
rect 552590 800 553618 856
rect 553786 800 554722 856
rect 554890 800 555918 856
rect 556086 800 557114 856
rect 557282 800 558310 856
rect 558478 800 559414 856
rect 559582 800 560610 856
rect 560778 800 561806 856
rect 561974 800 562910 856
rect 563078 800 564106 856
rect 564274 800 565302 856
rect 565470 800 566406 856
rect 566574 800 567602 856
rect 567770 800 568798 856
rect 568966 800 569902 856
rect 570070 800 571098 856
rect 571266 800 572294 856
rect 572462 800 573398 856
rect 573566 800 574594 856
rect 574762 800 575790 856
rect 575958 800 576894 856
rect 577062 800 577742 856
<< metal3 >>
rect 0 572568 800 572688
rect 579200 557064 580000 557184
rect 0 518032 800 518152
rect 579200 471384 580000 471504
rect 0 463496 800 463616
rect 0 408960 800 409080
rect 579200 385704 580000 385824
rect 0 354424 800 354544
rect 0 299888 800 300008
rect 579200 299888 580000 300008
rect 0 245352 800 245472
rect 579200 214208 580000 214328
rect 0 190816 800 190936
rect 0 136280 800 136400
rect 579200 128528 580000 128648
rect 0 81744 800 81864
rect 579200 42848 580000 42968
rect 0 27208 800 27328
<< obsm3 >>
rect 565 572768 579200 597345
rect 880 572488 579200 572768
rect 565 557264 579200 572488
rect 565 556984 579120 557264
rect 565 518232 579200 556984
rect 880 517952 579200 518232
rect 565 471584 579200 517952
rect 565 471304 579120 471584
rect 565 463696 579200 471304
rect 880 463416 579200 463696
rect 565 409160 579200 463416
rect 880 408880 579200 409160
rect 565 385904 579200 408880
rect 565 385624 579120 385904
rect 565 354624 579200 385624
rect 880 354344 579200 354624
rect 565 300088 579200 354344
rect 880 299808 579120 300088
rect 565 245552 579200 299808
rect 880 245272 579200 245552
rect 565 214408 579200 245272
rect 565 214128 579120 214408
rect 565 191016 579200 214128
rect 880 190736 579200 191016
rect 565 136480 579200 190736
rect 880 136200 579200 136480
rect 565 128728 579200 136200
rect 565 128448 579120 128728
rect 565 81944 579200 128448
rect 880 81664 579200 81944
rect 565 43048 579200 81664
rect 565 42768 579120 43048
rect 565 27408 579200 42768
rect 880 27128 579200 27408
rect 565 2143 579200 27128
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
rect 50288 2128 50608 597360
rect 65648 2128 65968 597360
rect 81008 2128 81328 597360
rect 96368 2128 96688 597360
rect 111728 2128 112048 597360
rect 127088 2128 127408 597360
rect 142448 2128 142768 597360
rect 157808 2128 158128 597360
rect 173168 2128 173488 597360
rect 188528 2128 188848 597360
rect 203888 2128 204208 597360
rect 219248 2128 219568 597360
rect 234608 2128 234928 597360
rect 249968 2128 250288 597360
rect 265328 2128 265648 597360
rect 280688 2128 281008 597360
rect 296048 2128 296368 597360
rect 311408 2128 311728 597360
rect 326768 2128 327088 597360
rect 342128 2128 342448 597360
rect 357488 2128 357808 597360
rect 372848 2128 373168 597360
rect 388208 2128 388528 597360
rect 403568 2128 403888 597360
rect 418928 2128 419248 597360
rect 434288 2128 434608 597360
rect 449648 2128 449968 597360
rect 465008 2128 465328 597360
rect 480368 2128 480688 597360
rect 495728 2128 496048 597360
rect 511088 2128 511408 597360
rect 526448 2128 526768 597360
rect 541808 2128 542128 597360
rect 557168 2128 557488 597360
rect 572528 2128 572848 597360
<< obsm4 >>
rect 48267 3435 50208 13973
rect 50688 3435 52381 13973
<< labels >>
rlabel metal2 s 572350 0 572406 800 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 0 190816 800 190936 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 579200 299888 580000 300008 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 0 245352 800 245472 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 0 299888 800 300008 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 567934 599200 567990 600000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 575846 0 575902 800 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 576950 0 577006 800 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 578146 0 578202 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 354424 800 354544 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 572718 599200 572774 600000 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 0 27208 800 27328 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 579200 385704 580000 385824 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 408960 800 409080 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 579200 471384 580000 471504 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 463496 800 463616 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 518032 800 518152 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 579200 557064 580000 557184 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 572568 800 572688 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal2 s 579342 0 579398 800 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 577502 599200 577558 600000 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 579200 128528 580000 128648 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal2 s 573454 0 573510 800 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal2 s 558366 599200 558422 600000 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 0 81744 800 81864 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal2 s 563150 599200 563206 600000 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 579200 214208 580000 214328 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal3 s 0 136280 800 136400 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 574650 0 574706 800 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 2410 599200 2466 600000 6 io_in[0]
port 30 nsew signal input
rlabel metal2 s 146114 599200 146170 600000 6 io_in[10]
port 31 nsew signal input
rlabel metal2 s 160558 599200 160614 600000 6 io_in[11]
port 32 nsew signal input
rlabel metal2 s 174910 599200 174966 600000 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 189262 599200 189318 600000 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 203706 599200 203762 600000 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 218058 599200 218114 600000 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 232410 599200 232466 600000 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 246854 599200 246910 600000 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 261206 599200 261262 600000 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 275558 599200 275614 600000 6 io_in[19]
port 40 nsew signal input
rlabel metal2 s 16762 599200 16818 600000 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 289910 599200 289966 600000 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 304354 599200 304410 600000 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 318706 599200 318762 600000 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 333058 599200 333114 600000 6 io_in[23]
port 45 nsew signal input
rlabel metal2 s 347502 599200 347558 600000 6 io_in[24]
port 46 nsew signal input
rlabel metal2 s 361854 599200 361910 600000 6 io_in[25]
port 47 nsew signal input
rlabel metal2 s 376206 599200 376262 600000 6 io_in[26]
port 48 nsew signal input
rlabel metal2 s 390650 599200 390706 600000 6 io_in[27]
port 49 nsew signal input
rlabel metal2 s 405002 599200 405058 600000 6 io_in[28]
port 50 nsew signal input
rlabel metal2 s 419354 599200 419410 600000 6 io_in[29]
port 51 nsew signal input
rlabel metal2 s 31114 599200 31170 600000 6 io_in[2]
port 52 nsew signal input
rlabel metal2 s 433706 599200 433762 600000 6 io_in[30]
port 53 nsew signal input
rlabel metal2 s 448150 599200 448206 600000 6 io_in[31]
port 54 nsew signal input
rlabel metal2 s 462502 599200 462558 600000 6 io_in[32]
port 55 nsew signal input
rlabel metal2 s 476854 599200 476910 600000 6 io_in[33]
port 56 nsew signal input
rlabel metal2 s 491298 599200 491354 600000 6 io_in[34]
port 57 nsew signal input
rlabel metal2 s 505650 599200 505706 600000 6 io_in[35]
port 58 nsew signal input
rlabel metal2 s 520002 599200 520058 600000 6 io_in[36]
port 59 nsew signal input
rlabel metal2 s 534446 599200 534502 600000 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 45466 599200 45522 600000 6 io_in[3]
port 61 nsew signal input
rlabel metal2 s 59910 599200 59966 600000 6 io_in[4]
port 62 nsew signal input
rlabel metal2 s 74262 599200 74318 600000 6 io_in[5]
port 63 nsew signal input
rlabel metal2 s 88614 599200 88670 600000 6 io_in[6]
port 64 nsew signal input
rlabel metal2 s 103058 599200 103114 600000 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 117410 599200 117466 600000 6 io_in[8]
port 66 nsew signal input
rlabel metal2 s 131762 599200 131818 600000 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 7194 599200 7250 600000 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 150990 599200 151046 600000 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 165342 599200 165398 600000 6 io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 179694 599200 179750 600000 6 io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 194046 599200 194102 600000 6 io_oeb[13]
port 72 nsew signal output
rlabel metal2 s 208490 599200 208546 600000 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 222842 599200 222898 600000 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 237194 599200 237250 600000 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 251638 599200 251694 600000 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 265990 599200 266046 600000 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 280342 599200 280398 600000 6 io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 21546 599200 21602 600000 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 294786 599200 294842 600000 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 309138 599200 309194 600000 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 323490 599200 323546 600000 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 337842 599200 337898 600000 6 io_oeb[23]
port 83 nsew signal output
rlabel metal2 s 352286 599200 352342 600000 6 io_oeb[24]
port 84 nsew signal output
rlabel metal2 s 366638 599200 366694 600000 6 io_oeb[25]
port 85 nsew signal output
rlabel metal2 s 380990 599200 381046 600000 6 io_oeb[26]
port 86 nsew signal output
rlabel metal2 s 395434 599200 395490 600000 6 io_oeb[27]
port 87 nsew signal output
rlabel metal2 s 409786 599200 409842 600000 6 io_oeb[28]
port 88 nsew signal output
rlabel metal2 s 424138 599200 424194 600000 6 io_oeb[29]
port 89 nsew signal output
rlabel metal2 s 35898 599200 35954 600000 6 io_oeb[2]
port 90 nsew signal output
rlabel metal2 s 438582 599200 438638 600000 6 io_oeb[30]
port 91 nsew signal output
rlabel metal2 s 452934 599200 452990 600000 6 io_oeb[31]
port 92 nsew signal output
rlabel metal2 s 467286 599200 467342 600000 6 io_oeb[32]
port 93 nsew signal output
rlabel metal2 s 481638 599200 481694 600000 6 io_oeb[33]
port 94 nsew signal output
rlabel metal2 s 496082 599200 496138 600000 6 io_oeb[34]
port 95 nsew signal output
rlabel metal2 s 510434 599200 510490 600000 6 io_oeb[35]
port 96 nsew signal output
rlabel metal2 s 524786 599200 524842 600000 6 io_oeb[36]
port 97 nsew signal output
rlabel metal2 s 539230 599200 539286 600000 6 io_oeb[37]
port 98 nsew signal output
rlabel metal2 s 50250 599200 50306 600000 6 io_oeb[3]
port 99 nsew signal output
rlabel metal2 s 64694 599200 64750 600000 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 79046 599200 79102 600000 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 93398 599200 93454 600000 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 107842 599200 107898 600000 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 122194 599200 122250 600000 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 136546 599200 136602 600000 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 11978 599200 12034 600000 6 io_out[0]
port 106 nsew signal output
rlabel metal2 s 155774 599200 155830 600000 6 io_out[10]
port 107 nsew signal output
rlabel metal2 s 170126 599200 170182 600000 6 io_out[11]
port 108 nsew signal output
rlabel metal2 s 184478 599200 184534 600000 6 io_out[12]
port 109 nsew signal output
rlabel metal2 s 198922 599200 198978 600000 6 io_out[13]
port 110 nsew signal output
rlabel metal2 s 213274 599200 213330 600000 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 227626 599200 227682 600000 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 241978 599200 242034 600000 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 256422 599200 256478 600000 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 270774 599200 270830 600000 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 285126 599200 285182 600000 6 io_out[19]
port 116 nsew signal output
rlabel metal2 s 26330 599200 26386 600000 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 299570 599200 299626 600000 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 313922 599200 313978 600000 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 328274 599200 328330 600000 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 342718 599200 342774 600000 6 io_out[23]
port 121 nsew signal output
rlabel metal2 s 357070 599200 357126 600000 6 io_out[24]
port 122 nsew signal output
rlabel metal2 s 371422 599200 371478 600000 6 io_out[25]
port 123 nsew signal output
rlabel metal2 s 385774 599200 385830 600000 6 io_out[26]
port 124 nsew signal output
rlabel metal2 s 400218 599200 400274 600000 6 io_out[27]
port 125 nsew signal output
rlabel metal2 s 414570 599200 414626 600000 6 io_out[28]
port 126 nsew signal output
rlabel metal2 s 428922 599200 428978 600000 6 io_out[29]
port 127 nsew signal output
rlabel metal2 s 40682 599200 40738 600000 6 io_out[2]
port 128 nsew signal output
rlabel metal2 s 443366 599200 443422 600000 6 io_out[30]
port 129 nsew signal output
rlabel metal2 s 457718 599200 457774 600000 6 io_out[31]
port 130 nsew signal output
rlabel metal2 s 472070 599200 472126 600000 6 io_out[32]
port 131 nsew signal output
rlabel metal2 s 486514 599200 486570 600000 6 io_out[33]
port 132 nsew signal output
rlabel metal2 s 500866 599200 500922 600000 6 io_out[34]
port 133 nsew signal output
rlabel metal2 s 515218 599200 515274 600000 6 io_out[35]
port 134 nsew signal output
rlabel metal2 s 529570 599200 529626 600000 6 io_out[36]
port 135 nsew signal output
rlabel metal2 s 544014 599200 544070 600000 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 55126 599200 55182 600000 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 69478 599200 69534 600000 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 83830 599200 83886 600000 6 io_out[5]
port 139 nsew signal output
rlabel metal2 s 98182 599200 98238 600000 6 io_out[6]
port 140 nsew signal output
rlabel metal2 s 112626 599200 112682 600000 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 126978 599200 127034 600000 6 io_out[8]
port 142 nsew signal output
rlabel metal2 s 141330 599200 141386 600000 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 474278 0 474334 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 477774 0 477830 800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 481270 0 481326 800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 484766 0 484822 800 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 488262 0 488318 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 491850 0 491906 800 6 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 495346 0 495402 800 6 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 498842 0 498898 800 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 502338 0 502394 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 505834 0 505890 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 509330 0 509386 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 512826 0 512882 800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 516322 0 516378 800 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 519818 0 519874 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 523314 0 523370 800 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 526810 0 526866 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 530306 0 530362 800 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 533802 0 533858 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 537298 0 537354 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 540794 0 540850 800 6 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 544290 0 544346 800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 547786 0 547842 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 551282 0 551338 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 554778 0 554834 800 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 558366 0 558422 800 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 561862 0 561918 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 565358 0 565414 800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 568854 0 568910 800 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 166262 0 166318 800 6 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 180246 0 180302 800 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 187238 0 187294 800 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 190734 0 190790 800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 194230 0 194286 800 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 201222 0 201278 800 6 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 208214 0 208270 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 211710 0 211766 800 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 215206 0 215262 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 225786 0 225842 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 229282 0 229338 800 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 236274 0 236330 800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 239770 0 239826 800 6 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 243266 0 243322 800 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 246762 0 246818 800 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 250258 0 250314 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 253754 0 253810 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 260746 0 260802 800 6 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 264242 0 264298 800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 267738 0 267794 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 271234 0 271290 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 274730 0 274786 800 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 278226 0 278282 800 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 281722 0 281778 800 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 285218 0 285274 800 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 288714 0 288770 800 6 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 292302 0 292358 800 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 295798 0 295854 800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 299294 0 299350 800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 306286 0 306342 800 6 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 309782 0 309838 800 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 313278 0 313334 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 316774 0 316830 800 6 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 320270 0 320326 800 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 323766 0 323822 800 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 327262 0 327318 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 330758 0 330814 800 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 334254 0 334310 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 337750 0 337806 800 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 341246 0 341302 800 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 344742 0 344798 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 348238 0 348294 800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 351734 0 351790 800 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 355230 0 355286 800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 358818 0 358874 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 362314 0 362370 800 6 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 365810 0 365866 800 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 369306 0 369362 800 6 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 372802 0 372858 800 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 376298 0 376354 800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 379794 0 379850 800 6 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 383290 0 383346 800 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 386786 0 386842 800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 390282 0 390338 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 393778 0 393834 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 397274 0 397330 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 400770 0 400826 800 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 404266 0 404322 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 407762 0 407818 800 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 411258 0 411314 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 414754 0 414810 800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 418250 0 418306 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 421746 0 421802 800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 425334 0 425390 800 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 428830 0 428886 800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 432326 0 432382 800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 435822 0 435878 800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 439318 0 439374 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 442814 0 442870 800 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 446310 0 446366 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 449806 0 449862 800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 453302 0 453358 800 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 456798 0 456854 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 460294 0 460350 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 463790 0 463846 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 467286 0 467342 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 470782 0 470838 800 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 475474 0 475530 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 478970 0 479026 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 482466 0 482522 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 485962 0 486018 800 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 489458 0 489514 800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 492954 0 493010 800 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 496450 0 496506 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 499946 0 500002 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 503442 0 503498 800 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 506938 0 506994 800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 510434 0 510490 800 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 514022 0 514078 800 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 517518 0 517574 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 521014 0 521070 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 524510 0 524566 800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 528006 0 528062 800 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 531502 0 531558 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 534998 0 535054 800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 538494 0 538550 800 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 541990 0 542046 800 6 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 545486 0 545542 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 548982 0 549038 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 552478 0 552534 800 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 555974 0 556030 800 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 559470 0 559526 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 562966 0 563022 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 566462 0 566518 800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 569958 0 570014 800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 167366 0 167422 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 170862 0 170918 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 177854 0 177910 800 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 181442 0 181498 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 184938 0 184994 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 188434 0 188490 800 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 191930 0 191986 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 128910 0 128966 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 195426 0 195482 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 198922 0 198978 800 6 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 202418 0 202474 800 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 205914 0 205970 800 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 209410 0 209466 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 212906 0 212962 800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 216402 0 216458 800 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 219898 0 219954 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 223394 0 223450 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 226890 0 226946 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 132406 0 132462 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 230386 0 230442 800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 233882 0 233938 800 6 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 237378 0 237434 800 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 240874 0 240930 800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 244370 0 244426 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 247958 0 248014 800 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 251454 0 251510 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 254950 0 255006 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 258446 0 258502 800 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 261942 0 261998 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 265438 0 265494 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 268934 0 268990 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 272430 0 272486 800 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 275926 0 275982 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 279422 0 279478 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 282918 0 282974 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 286414 0 286470 800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 289910 0 289966 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 293406 0 293462 800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 296902 0 296958 800 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 300398 0 300454 800 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 303894 0 303950 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 307390 0 307446 800 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 310886 0 310942 800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 314474 0 314530 800 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 317970 0 318026 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 321466 0 321522 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 324962 0 325018 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 328458 0 328514 800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 331954 0 332010 800 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 335450 0 335506 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 338946 0 339002 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 342442 0 342498 800 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 345938 0 345994 800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 349434 0 349490 800 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 352930 0 352986 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 356426 0 356482 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 359922 0 359978 800 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 363418 0 363474 800 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 366914 0 366970 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 146390 0 146446 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 370410 0 370466 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 373906 0 373962 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 377402 0 377458 800 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 380990 0 381046 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 384486 0 384542 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 387982 0 388038 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 391478 0 391534 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 394974 0 395030 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 398470 0 398526 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 401966 0 402022 800 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 149886 0 149942 800 6 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 405462 0 405518 800 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 408958 0 409014 800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 412454 0 412510 800 6 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 415950 0 416006 800 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 419446 0 419502 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 422942 0 422998 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 426438 0 426494 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 429934 0 429990 800 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 433430 0 433486 800 6 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 436926 0 436982 800 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 153382 0 153438 800 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 440422 0 440478 800 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 443918 0 443974 800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 447506 0 447562 800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 451002 0 451058 800 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 454498 0 454554 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 457994 0 458050 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 461490 0 461546 800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 464986 0 465042 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 468482 0 468538 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 471978 0 472034 800 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 156878 0 156934 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 126518 0 126574 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 476670 0 476726 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 480166 0 480222 800 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 483662 0 483718 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 487158 0 487214 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 490654 0 490710 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 494150 0 494206 800 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 497646 0 497702 800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 501142 0 501198 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 504638 0 504694 800 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 508134 0 508190 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 511630 0 511686 800 6 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 515126 0 515182 800 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 518622 0 518678 800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 522118 0 522174 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 525614 0 525670 800 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 529110 0 529166 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 532606 0 532662 800 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 536194 0 536250 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 539690 0 539746 800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 543186 0 543242 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 546682 0 546738 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 550178 0 550234 800 6 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 553674 0 553730 800 6 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 557170 0 557226 800 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 560666 0 560722 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 564162 0 564218 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 567658 0 567714 800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 571154 0 571210 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 182546 0 182602 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 186042 0 186098 800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 200026 0 200082 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 203614 0 203670 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 207110 0 207166 800 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 210606 0 210662 800 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 214102 0 214158 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 217598 0 217654 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 221094 0 221150 800 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 224590 0 224646 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 228086 0 228142 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 231582 0 231638 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 238574 0 238630 800 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 242070 0 242126 800 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 249062 0 249118 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 252558 0 252614 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 256054 0 256110 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 266542 0 266598 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 270130 0 270186 800 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 273626 0 273682 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 277122 0 277178 800 6 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 280618 0 280674 800 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 284114 0 284170 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 287610 0 287666 800 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 291106 0 291162 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 294602 0 294658 800 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 298098 0 298154 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 301594 0 301650 800 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 305090 0 305146 800 6 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 308586 0 308642 800 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 312082 0 312138 800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 315578 0 315634 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 319074 0 319130 800 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 322570 0 322626 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 326066 0 326122 800 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 329562 0 329618 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 333058 0 333114 800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 336646 0 336702 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 340142 0 340198 800 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 343638 0 343694 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 347134 0 347190 800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 350630 0 350686 800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 354126 0 354182 800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 357622 0 357678 800 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 361118 0 361174 800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 364614 0 364670 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 368110 0 368166 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 371606 0 371662 800 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 375102 0 375158 800 6 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 378598 0 378654 800 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 382094 0 382150 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 385590 0 385646 800 6 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 389086 0 389142 800 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 392582 0 392638 800 6 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 396078 0 396134 800 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 399574 0 399630 800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 403162 0 403218 800 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 406658 0 406714 800 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 410154 0 410210 800 6 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 413650 0 413706 800 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 417146 0 417202 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 420642 0 420698 800 6 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 424138 0 424194 800 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 427634 0 427690 800 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 431130 0 431186 800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 434626 0 434682 800 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 438122 0 438178 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 441618 0 441674 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 445114 0 445170 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 448610 0 448666 800 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 452106 0 452162 800 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 455602 0 455658 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 459098 0 459154 800 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 462594 0 462650 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 466090 0 466146 800 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 469678 0 469734 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 473174 0 473230 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_oenb[9]
port 527 nsew signal input
rlabel metal3 s 579200 42848 580000 42968 6 user_irq[0]
port 528 nsew signal output
rlabel metal2 s 548798 599200 548854 600000 6 user_irq[1]
port 529 nsew signal output
rlabel metal2 s 553582 599200 553638 600000 6 user_irq[2]
port 530 nsew signal output
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 65648 2128 65968 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 96368 2128 96688 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 127088 2128 127408 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 157808 2128 158128 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 188528 2128 188848 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 219248 2128 219568 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 249968 2128 250288 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 280688 2128 281008 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 311408 2128 311728 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 342128 2128 342448 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 372848 2128 373168 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 403568 2128 403888 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 434288 2128 434608 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 465008 2128 465328 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 495728 2128 496048 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 526448 2128 526768 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 557168 2128 557488 597360 6 vccd1
port 531 nsew power input
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 50288 2128 50608 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 81008 2128 81328 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 111728 2128 112048 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 142448 2128 142768 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 173168 2128 173488 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 203888 2128 204208 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 234608 2128 234928 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 265328 2128 265648 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 296048 2128 296368 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 326768 2128 327088 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 357488 2128 357808 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 388208 2128 388528 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 418928 2128 419248 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 449648 2128 449968 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 480368 2128 480688 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 511088 2128 511408 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 541808 2128 542128 597360 6 vssd1
port 532 nsew ground input
rlabel metal4 s 572528 2128 572848 597360 6 vssd1
port 532 nsew ground input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 533 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 534 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_ack_o
port 535 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[0]
port 536 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 wbs_adr_i[10]
port 537 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wbs_adr_i[11]
port 538 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 wbs_adr_i[12]
port 539 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wbs_adr_i[13]
port 540 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wbs_adr_i[14]
port 541 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 wbs_adr_i[15]
port 542 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 wbs_adr_i[16]
port 543 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 wbs_adr_i[17]
port 544 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 wbs_adr_i[18]
port 545 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 wbs_adr_i[19]
port 546 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_adr_i[1]
port 547 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 wbs_adr_i[20]
port 548 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 wbs_adr_i[21]
port 549 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 wbs_adr_i[22]
port 550 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 wbs_adr_i[23]
port 551 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 wbs_adr_i[24]
port 552 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 wbs_adr_i[25]
port 553 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 wbs_adr_i[26]
port 554 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 wbs_adr_i[27]
port 555 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 wbs_adr_i[28]
port 556 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 wbs_adr_i[29]
port 557 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[2]
port 558 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 wbs_adr_i[30]
port 559 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 wbs_adr_i[31]
port 560 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[3]
port 561 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[4]
port 562 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[5]
port 563 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_adr_i[6]
port 564 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_adr_i[7]
port 565 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_adr_i[8]
port 566 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_adr_i[9]
port 567 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_cyc_i
port 568 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_i[0]
port 569 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 wbs_dat_i[10]
port 570 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 wbs_dat_i[11]
port 571 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_dat_i[12]
port 572 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_i[13]
port 573 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 wbs_dat_i[14]
port 574 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 wbs_dat_i[15]
port 575 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 wbs_dat_i[16]
port 576 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 wbs_dat_i[17]
port 577 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 wbs_dat_i[18]
port 578 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 wbs_dat_i[19]
port 579 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_i[1]
port 580 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 wbs_dat_i[20]
port 581 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 wbs_dat_i[21]
port 582 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 wbs_dat_i[22]
port 583 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 wbs_dat_i[23]
port 584 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 wbs_dat_i[24]
port 585 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 wbs_dat_i[25]
port 586 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 wbs_dat_i[26]
port 587 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 wbs_dat_i[27]
port 588 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 wbs_dat_i[28]
port 589 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 wbs_dat_i[29]
port 590 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[2]
port 591 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 wbs_dat_i[30]
port 592 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 wbs_dat_i[31]
port 593 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_i[3]
port 594 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_i[4]
port 595 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_i[5]
port 596 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_i[6]
port 597 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[7]
port 598 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_dat_i[8]
port 599 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_i[9]
port 600 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[0]
port 601 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 wbs_dat_o[10]
port 602 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_o[11]
port 603 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 wbs_dat_o[12]
port 604 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 wbs_dat_o[13]
port 605 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 wbs_dat_o[14]
port 606 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 wbs_dat_o[15]
port 607 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 wbs_dat_o[16]
port 608 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 wbs_dat_o[17]
port 609 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 wbs_dat_o[18]
port 610 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 wbs_dat_o[19]
port 611 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[1]
port 612 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 wbs_dat_o[20]
port 613 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 wbs_dat_o[21]
port 614 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 wbs_dat_o[22]
port 615 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 wbs_dat_o[23]
port 616 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 wbs_dat_o[24]
port 617 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 wbs_dat_o[25]
port 618 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 wbs_dat_o[26]
port 619 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 wbs_dat_o[27]
port 620 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 wbs_dat_o[28]
port 621 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 wbs_dat_o[29]
port 622 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_o[2]
port 623 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 wbs_dat_o[30]
port 624 nsew signal output
rlabel metal2 s 123022 0 123078 800 6 wbs_dat_o[31]
port 625 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_o[3]
port 626 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_o[4]
port 627 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[5]
port 628 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_o[6]
port 629 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_o[7]
port 630 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_o[8]
port 631 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_o[9]
port 632 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_sel_i[0]
port 633 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_sel_i[1]
port 634 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_sel_i[2]
port 635 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_sel_i[3]
port 636 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_stb_i
port 637 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_we_i
port 638 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 580000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 90222184
string GDS_FILE /home/ren/Projects/caravel_tutorial/caravel_example/openlane/NNgen/runs/NNgen/results/finishing/basic.magic.gds
string GDS_START 190330
<< end >>

